module dm_4k(addr, din, MemWrite, clk, dout);
    input [11:2] addr;           // address bus
    input [31:0] din;            // 32-bit input data
    input MemWrite;                    // memory write enable
    input clk;                   // clock
    output reg [31:0] dout;      // 32-bit memory output

    reg [31:0] dm[1023:0];

    integer i;
    initial begin
      for (i = 0; i < 1024 ; i = i + 1) begin
          dm[i] <= 0;
      end
    end

    always @(posedge clk) begin
        if(MemWrite) begin
            dm[addr] <= din;
        end
        else dout <= dm[addr];
    end
endmodule
