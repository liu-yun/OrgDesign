module im_4k(addr, dout);
    input [11:2] addr;  // address bus
    output [31:0] dout; // 32-bit memory output

    reg [31:0] im[1023:0];
    integer i;

    initial begin
      for (i = 0; i < 1024 ; i = i + 1) begin
          im[i] = 0;
      end
      $readmemh("code.txt", im);
    end
    
    assign dout = im[addr];
endmodule
